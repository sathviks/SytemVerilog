/*  Modport    */


/*

=>  The Modport groups and specifies the port directions to the wires/signals declared within the interface.
     modports are declared inside the interface with the keyword modport.


     It help us to prevent wireing errors





Example :

    Monitor should be never be driving input signals similarly driver should not be driving output signals


 //modport delcaration
  modport driver  (input a, output b);
  modport monitor (input a, input  b);

*/


interface add_if;
  logic [3:0] a;
  logic [3:0] b;
  logic [4:0] sum;
  logic clk;
  
  modport DRV (output a,b, input sum,clk);
  modport MON (output sum,clk, input a,b);
 
  
endinterface
 
 
class driver;
  
  virtual add_if.DRV aif; //declaration
  
  task run();
    forever begin
      @(posedge aif.clk);  
      aif.a <= 2;
      aif.b <= 3;
      $display("[DRV] : Interface Trigger");
    end
  endtask
  
  
endclass
 
 
 
module tb;
  
 add_if aif();
  driver drv;
  
  add dut (aif.a, aif.b, aif.sum, aif.clk );
 
 
  initial begin
    aif.clk <= 0;
  end
  
  always #10 aif.clk <= ~aif.clk;
 
   initial begin
     drv = new();
     drv.aif = aif;
     drv.run();
     
   end
  
  initial begin
    $dumpfile("dump.vcd"); 
    $dumpvars;  
    #100;
    $finish();
  end
  
endmodule